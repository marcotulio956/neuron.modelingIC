module izhikevich_neuron #() ();

endmodule